FDISK

FDISK �r ett grundverktyg f�r att ta bort och skapa partitioner p� h�rddiskar
