Begin3
Language:    SV, 850, Swedish
Title:       Free FDISK
Description: Verktyg f�r fixa diskar - skapa partitioner.
Keywords:    fdisk, formatera, h�rddisk, partition, fat16, fat32, partition, mbr
End
